
`include "parameters.sv"  
`include "ALU.sv"
`include "regfile.sv"
`include "mux.sv"
`include "decode.sv"
`include "instruction_memory.sv"
`include "data_memory.sv"
`include "fsm_control.sv"
`include "datapath.sv"
`include "cpu.sv"


